`define INT 8'hc0 // format B
`define IRET 8'hc0 // format B
`define IRES 8'hc0 // format B
`define WAIT 8'hc0 // format B
`define LCTRL 8'ha0 // format F
`define SCTRL 8'ha1 // format F
`define FLAG 8'h80 // format I
`define ADDIP 8'h81 // format I
`define JAL 8'h82 // format I
`define JALR 8'h83 // format I
`define RET 8'h84 // format I
`define RETR 8'h85 // format I
`define BRA 8'hc1 // format B
`define BEQ 8'hc1 // format B
`define BEZ 8'hc1 // format B
`define BLT 8'hc1 // format B
`define BLE 8'hc1 // format B
`define BLTU 8'hc1 // format B
`define BLEU 8'hc1 // format B
`define BNE 8'hc1 // format B
`define BNZ 8'hc1 // format B
`define BGE 8'hc1 // format B
`define BGT 8'hc1 // format B
`define BGEU 8'hc1 // format B
`define BGTU 8'hc1 // format B
`define PUSH 8'h86 // format I
`define POP 8'h87 // format I
`define ENTER 8'h88 // format I
`define LEAVE 8'h89 // format I
`define CMP 8'h8a // format I
`define LLI 8'ha2 // format F
`define LLIP 8'ha2 // format F
`define LNI 8'he0 // format U
`define LTI 8'he1 // format U
`define LW 8'h20 // format E
`define LH 8'h21 // format E
`define LHS 8'h22 // format E
`define LQ 8'h23 // format E
`define LQS 8'h24 // format E
`define LB 8'h25 // format E
`define LBS 8'h26 // format E
`define SW 8'h27 // format E
`define SH 8'h28 // format E
`define SQ 8'h29 // format E
`define SB 8'h2a // format E
`define LLW 8'h3f // format E
`define LLH 8'h3f // format E
`define LLQ 8'h3f // format E
`define LLB 8'h3f // format E
`define SCW 8'h3f // format E
`define SCH 8'h3f // format E
`define SCQ 8'h3f // format E
`define SCB 8'h3f // format E
`define LFENCE 8'hc3 // format B
`define SFENCE 8'hc3 // format B
`define MFENCE 8'hc3 // format B
`define TFLUSHX 8'hc3 // format B
`define TFLUSH 8'hc3 // format B
`define ADDR 8'h40 // format R
`define ADDI 8'h8b // format I
`define IADC 8'h41 // format R
`define UADC 8'h41 // format R
`define SUBR 8'h42 // format R
`define SUBI 8'h8c // format I
`define ISBB 8'h43 // format R
`define USBB 8'h43 // format R
`define IMULR 8'h44 // format R
`define IMULH 8'h45 // format R
`define IMULI 8'h8c // format I
`define IDIVR 8'h46 // format R
`define IDIVI 8'h8e // format I
`define UMULR 8'h47 // format R
`define UMULH 8'h48 // format R
`define UMULI 8'h8f // format I
`define UDIVR 8'h49 // format R
`define UDIVI 8'h90 // format I
`define REMR 8'h4a // format R
`define REMI 8'h91 // format I
`define MODR 8'h4b // format R
`define MODI 8'h92 // format I
`define ANDR 8'h4c // format R
`define ANDI 8'h93 // format I
`define ORR 8'h4d // format R
`define ORI 8'h94 // format I
`define NORR 8'h4e // format R
`define NORI 8'h95 // format I
`define XORR 8'h4f // format R
`define XORI 8'h96 // format I
`define SHL 8'h50 // format R
`define ASR 8'h51 // format R
`define LSR 8'h52 // format R
`define FCMP 8'h2b // format E
`define FTO 8'h2c // format E
`define FFROM 8'h2d // format E
`define FNEG 8'h2e // format E
`define FABS 8'h2f // format E
`define FADD 8'h30 // format E
`define FSUB 8'h31 // format E
`define FMUL 8'h32 // format E
`define FDIV 8'h33 // format E
`define FMA 8'h34 // format E
`define FSQRT 8'h35 // format E
`define FMIN 8'h36 // format E
`define FMAX 8'h37 // format E
`define FRND 8'h38 // format E
`define FRNDA 8'h38 // format E
`define FTRUNC 8'h38 // format E
`define FCEIL 8'h38 // format E
`define FFLOOR 8'h38 // format E
`define FCNV 8'h39 // format E
`define FCLASS 8'h3a // format E
`define RORR 8'h53 // format R
`define RORI 8'h97 // format I
`define ROLR 8'h54 // format R
`define ROLI 8'h98 // format I
`define CSET 8'h55 // format R
`define CLZ 8'h56 // format R
`define CTZ 8'h57 // format R
`define EXT 8'h58 // format R
`define DEP 8'h59 // format R
`define ZIP 8'h99 // format I
`define REV 8'h9a // format I
`define ANDN 8'h5a // format R
`define ORN 8'h5b // format R
`define XORN 8'h5c // format R
